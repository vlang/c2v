module main

const builtins = ''
