[translated]
module main

fn main()  {
        pointers := [8]&void{}
        return
}