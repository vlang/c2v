[translated]
module main


[typedef]
struct C.FILE {}


// vstart

fn main()  {
	a := 0
	if (a = C.puts(c'Hello World')) {
		C.puts(c'noes')
	}
	if (a = C.puts(c'Hello World')) != 0 {
		C.puts(c'noes')
	}
	cacatua := 0
	if (cacatua = C.puts(c'Hello World')) {
		C.puts(c'noes')
	}
}

